`include "mycpu_top.h"

module id_stage(
    input clk,
    input reset,

    // pipeline control
    output id_allow_in,
    input  if_to_id_valid,
    input  exe_allow_in,
    output id_to_exe_valid,

    // bus from if
    input [`IF_TO_ID_BUS_WIDTH-1:0] if_to_id_bus,

    // bus to exe
    output [`ID_TO_EXE_BUS_WIDTH-1:0] id_to_exe_bus,

    // buses from downstream stages (hazard detect)
    input [`EXE_TO_ID_BUS_WIDTH-1:0] exe_to_id_bus,
    input [`MEM_TO_ID_BUS_WIDTH-1:0] mem_to_id_bus,

    // bus to if (for branch)
    output [`ID_TO_IF_BUS_WIDTH-1:0] id_to_if_bus,

    // bus from wb (for regfile)
    input [`WB_TO_ID_BUS_WIDTH-1:0] wb_to_id_bus,

    // branch predictor update interface
    output        upd_en,
    output [31:0] upd_inst_addr,
    output        upd_br_inst,
    output        upd_cond_br_inst,
    output        upd_br_taken,
    output [31:0] upd_br_target
);

    // pipeline registers
    reg [`IF_TO_ID_BUS_WIDTH-1:0] id_reg;
    wire [31:0] id_pc;
    wire [31:0] id_inst;
    wire        id_pred_br_taken_X;
    reg         id_pred_br_taken;
    assign {id_pred_br_taken_X, id_pc, id_inst} = id_reg;
    // assign id_pred_br_taken = if_to_id_bus[64];
    

    // input bus from WB
    wire        wb_valid;
    wire        wb_rf_we_raw;
    wire [4:0]  wb_rf_waddr;
    wire [31:0] wb_rf_wdata;
    assign {wb_valid, wb_rf_we_raw, wb_rf_waddr, wb_rf_wdata} = wb_to_id_bus;

    // Hazard Detect
    wire        exe_valid;
    wire        exe_rf_we_raw;
    wire [4:0]  exe_rf_waddr;
    wire [31:0] exe_rf_wdata;
    wire        exe_is_load;
    assign {exe_valid, exe_rf_we_raw, exe_rf_waddr, exe_rf_wdata, exe_is_load} = exe_to_id_bus;
    
    wire        mem_valid;
    wire        mem_rf_we_raw;
    wire [4:0]  mem_rf_waddr;
    wire [31:0] mem_rf_wdata;
    wire        mem_is_load; // NEW: 从 MEM 段获取是否为 Load 指令
    assign {mem_valid, mem_rf_we_raw, mem_rf_waddr, mem_rf_wdata, mem_is_load} = mem_to_id_bus;

    wire wb_rf_we = wb_valid && wb_rf_we_raw;
    wire exe_rf_we = exe_valid && exe_rf_we_raw;
    wire mem_rf_we = mem_valid && mem_rf_we_raw;

    // output bus signals
    wire [31:0] rj_value;
    wire [31:0] rkd_value;
    wire [31:0] imm;
    wire [11:0] alu_op;
    wire        src1_is_pc;
    wire        src2_is_imm;
    wire        res_from_mem;
    wire        reg_we;
    wire        mem_en;
    wire [3:0]  mem_we;
    wire [4:0]  reg_waddr;
    wire [1:0]  data_sram_size; // New: 2'b00 Byte, 2'b10 Word

    assign id_to_exe_bus = {
        id_pc,       
        rj_value,    
        rkd_value,   
        imm,         
        alu_op,      
        src1_is_pc,  
        src2_is_imm, 
        res_from_mem,
        reg_we,      
        mem_en,      
        mem_we,      
        reg_waddr,
        data_sram_size // 传递给 EXE
    };

    // Branch bus
    wire        actual_br_taken;
    wire        br_cancel;
    reg         cancel_next;
    wire [31:0] br_target;
    wire [31:0] actual_br_target;
    assign id_to_if_bus = {actual_br_taken, actual_br_target};

    // Decoder Signals
    wire [5:0]  op_31_26;
    wire [3:0]  op_25_22;
    wire [1:0]  op_21_20;
    wire [4:0]  op_19_15;
    wire [4:0]  rd;
    wire [4:0]  rj;
    wire [4:0]  rk;
    wire [11:0] i12;
    wire [19:0] i20;
    wire [15:0] i16;
    wire [25:0] i26;

    assign op_31_26 = id_inst[31:26];
    assign op_25_22 = id_inst[25:22];
    assign op_21_20 = id_inst[21:20];
    assign op_19_15 = id_inst[19:15];
    assign rd   = id_inst[4:0];
    assign rj   = id_inst[9:5];
    assign rk   = id_inst[14:10];
    assign i12  = id_inst[21:10];
    assign i20  = id_inst[24:5];
    assign i16  = id_inst[25:10];
    assign i26  = {id_inst[9:0], id_inst[25:10]};

    wire [63:0] op_31_26_d;
    wire [15:0] op_25_22_d;
    wire [3:0]  op_21_20_d;
    wire [31:0] op_19_15_d;

    decoder_6_64 u_dec0 (.in(op_31_26), .out(op_31_26_d));
    decoder_4_16 u_dec1 (.in(op_25_22), .out(op_25_22_d));
    decoder_2_4  u_dec2 (.in(op_21_20), .out(op_21_20_d));
    decoder_5_32 u_dec3 (.in(op_19_15), .out(op_19_15_d));

    // Instruction Decode (Added New Instructions)
    wire inst_add_w     = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h00];
    wire inst_sub_w     = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h02];
    wire inst_slt       = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h04];
    wire inst_sltu      = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h05];
    wire inst_nor       = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h08];
    wire inst_and       = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h09];
    wire inst_or        = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h0a];
    wire inst_xor       = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h0b]; // NEW: XOR
    wire inst_mul       = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h18];
    wire inst_slli_w    = op_31_26_d[6'h00] & op_25_22_d[4'h1] & op_21_20_d[2'h0] & op_19_15_d[5'h01];
    wire inst_srli_w    = op_31_26_d[6'h00] & op_25_22_d[4'h1] & op_21_20_d[2'h0] & op_19_15_d[5'h09]; // NEW: SRLI.W
    wire inst_srai_w    = op_31_26_d[6'h00] & op_25_22_d[4'h1] & op_21_20_d[2'h0] & op_19_15_d[5'h11];
    wire inst_addi_w    = op_31_26_d[6'h00] & op_25_22_d[4'ha];
    wire inst_andi      = op_31_26_d[6'h00] & op_25_22_d[4'hd]; // NEW: ANDI
    wire inst_ori       = op_31_26_d[6'h00] & op_25_22_d[4'he];
    wire inst_pcaddu12i = op_31_26_d[6'h07] & ~id_inst[25];     // NEW: PCADDU12I
    wire inst_ld_b      = op_31_26_d[6'h0a] & op_25_22_d[4'h0]; // NEW: LD.B
    wire inst_ld_w      = op_31_26_d[6'h0a] & op_25_22_d[4'h2];
    wire inst_st_b      = op_31_26_d[6'h0a] & op_25_22_d[4'h4]; // NEW: ST.B
    wire inst_st_w      = op_31_26_d[6'h0a] & op_25_22_d[4'h6];
    wire inst_slti      = op_31_26_d[6'h00] & op_25_22_d[4'h8];
    wire inst_jirl      = op_31_26_d[6'h13];
    wire inst_b         = op_31_26_d[6'h14];
    wire inst_bl        = op_31_26_d[6'h15];
    wire inst_beq       = op_31_26_d[6'h16];
    wire inst_bne       = op_31_26_d[6'h17];                    // NEW: BNE
    wire inst_lu12i_w   = op_31_26_d[6'h05] & ~id_inst[25];

    // ALU Op Code Mapping
    assign alu_op[0]  = inst_add_w | inst_addi_w | inst_ld_w | inst_st_w | inst_jirl | inst_bl | inst_pcaddu12i | inst_ld_b | inst_st_b; // add
    assign alu_op[1]  = inst_sub_w; 
    assign alu_op[2]  = inst_slt | inst_slti;
    assign alu_op[3]  = inst_sltu;
    assign alu_op[4]  = inst_and | inst_andi;
    assign alu_op[5]  = inst_xor; // Replaced NOR with XOR
    assign alu_op[6]  = inst_or | inst_ori;
    assign alu_op[7]  = inst_mul;
    assign alu_op[8]  = inst_slli_w;
    assign alu_op[9]  = inst_srli_w;
    assign alu_op[10] = inst_srai_w;
    assign alu_op[11] = inst_lu12i_w;

    // Immediate generation
    wire need_ui5  = inst_slli_w | inst_srli_w | inst_srai_w;
    wire need_si12 = inst_addi_w | inst_ld_w | inst_st_w | inst_slti | inst_ld_b | inst_st_b;
    wire need_si16 = inst_jirl | inst_beq | inst_bne;
    wire need_si20 = inst_lu12i_w | inst_pcaddu12i;
    wire need_si26 = inst_b | inst_bl;
    wire src2_is_4 = inst_jirl | inst_bl;
    wire need_ui12 = inst_ori | inst_andi; // ANDI also uses Zero Extended imm

    assign imm = src2_is_4 ? 32'h4 :
                 need_si20 ? {i20[19:0], 12'b0} :
                 need_ui12 ? {20'b0, i12[11:0]} : // Zero Extend
                 {{20{i12[11]}}, i12[11:0]};      // Sign Extend

    // Operands Select
    assign src_reg_is_rd = inst_beq | inst_bne | inst_st_w | inst_st_b;
    assign src1_is_pc = inst_jirl | inst_bl | inst_pcaddu12i; // PCADDU12I uses PC

    assign src2_is_imm = inst_slli_w |
                     inst_srli_w |
                     inst_srai_w |
                     inst_addi_w |
                     inst_ld_w |
                     inst_ld_b |
                     inst_st_w |
                     inst_st_b |
                     inst_lu12i_w |
                     inst_pcaddu12i |
                     inst_jirl |
                     inst_bl |
                     inst_ori |
                     inst_andi |
                     inst_slti;

    assign res_from_mem = inst_ld_w | inst_ld_b;
    wire dst_is_r1 = inst_bl;
    assign reg_waddr = dst_is_r1 ? 5'd1 : rd;
    assign reg_we = (~inst_st_w & ~inst_st_b & ~inst_beq & ~inst_bne & ~inst_b) && |(reg_waddr);

    assign mem_en = inst_ld_w || inst_st_w || inst_ld_b || inst_st_b;
    // Note: For st.b, we still send 1111 to EXE, and EXE handles strobe based on address.
    assign mem_we = {4{inst_st_w | inst_st_b}}; 

    // 00: Byte, 01: Half, 10: Word
    assign data_sram_size = (inst_ld_b | inst_st_b) ? 2'b00 : 2'b10;

    // Regfile Read
    wire [4:0] rf_raddr1;
    wire [4:0] rf_raddr2;
    wire [31:0] rf_rdata1;
    wire [31:0] rf_rdata2;

    assign rf_raddr1 = rj;
    assign rf_raddr2 = src_reg_is_rd ? rd : rk;

    regfile u_regfile (
        .clk    (clk),
        .raddr1 (rf_raddr1),
        .rdata1 (rf_rdata1),
        .raddr2 (rf_raddr2),
        .rdata2 (rf_rdata2),
        .we     (wb_rf_we),
        .waddr  (wb_rf_waddr),
        .wdata  (wb_rf_wdata)
    );

    // Hazard Detection / Bypass (Standard)
    assign rj_value = 
        (exe_valid && exe_rf_we && (rf_raddr1 == exe_rf_waddr)) ? exe_rf_wdata :
        (mem_valid && mem_rf_we && (rf_raddr1 == mem_rf_waddr)) ? mem_rf_wdata :
        (wb_valid  && wb_rf_we  && (rf_raddr1 == wb_rf_waddr )) ? wb_rf_wdata  :
        rf_rdata1;
    assign rkd_value = 
        (exe_valid && exe_rf_we && (rf_raddr2 == exe_rf_waddr)) ? exe_rf_wdata :
        (mem_valid && mem_rf_we && (rf_raddr2 == mem_rf_waddr)) ? mem_rf_wdata :
        (wb_valid  && wb_rf_we  && (rf_raddr2 == wb_rf_waddr )) ? wb_rf_wdata  :
        rf_rdata2;

    wire rj_eq_rd = (rj_value == rkd_value);

    // Branch Logic
    wire br_taken;
    wire inst_is_br;
    wire inst_is_cond_br;
    wire [31:0] br_offs;
    wire [31:0] jirl_offs;

    assign br_offs = need_si26 ? {{4{i26[25]}}, i26[25:0], 2'b0} : {{14{i16[15]}}, i16[15:0], 2'b0};
    assign jirl_offs = {{14{i16[15]}}, i16[15:0], 2'b0};

    assign inst_is_br = inst_beq || inst_bne || inst_jirl || inst_bl || inst_b;
    assign inst_is_cond_br = inst_beq || inst_bne;

    assign br_taken = id_valid && ( inst_beq && rj_eq_rd
                    || inst_bne && !rj_eq_rd // BNE condition
                    || inst_jirl
                    || inst_bl
                    || inst_b
                    );

    assign br_target = ((inst_beq || inst_bne || inst_bl || inst_b) ? (id_pc + br_offs) :
                    /*inst_jirl*/ (rj_value + jirl_offs));
    
    assign actual_br_target = (br_taken && !id_pred_br_taken) ? br_target: (id_pc + 32'h4);

    wire br_mispred;
    assign br_mispred = id_valid && (br_taken != id_pred_br_taken);
    assign actual_br_taken = id_valid && id_allow_in && br_mispred; 
    assign br_cancel = actual_br_taken;

    // Ready/Valid logic
    reg  id_valid;
    wire id_ready_go;
    wire use_rf_rdata1 = id_valid && (
        inst_add_w   || inst_sub_w   || inst_slt   || inst_sltu ||
        inst_nor     || inst_and     || inst_or    || inst_xor || inst_mul ||
        inst_slli_w  || inst_srli_w  || inst_srai_w ||
        inst_addi_w  || inst_andi    || inst_ori   || inst_slti ||
        inst_ld_w    || inst_ld_b    || inst_st_w  || inst_st_b || 
        inst_jirl    || inst_beq     || inst_bne
    );
    wire use_rf_rdata2 = id_valid && (
        inst_add_w   || inst_sub_w   || inst_slt   || inst_sltu ||
        inst_nor     || inst_and     || inst_or    || inst_xor || inst_mul ||
        inst_st_w    || inst_st_b    || inst_beq   || inst_bne
    );
    
    // wire rf_rdata1_hazard = use_rf_rdata1 && (exe_valid && exe_is_load && exe_rf_we && (rf_raddr1 == exe_rf_waddr));
    // wire rf_rdata2_hazard = use_rf_rdata2 && (exe_valid && exe_is_load && exe_rf_we && (rf_raddr2 == exe_rf_waddr));
    // 检测 EXE 段的 Load 冲突
    // 检测 MEM 段的 Load 冲突
    wire rf_rdata1_hazard = use_rf_rdata1 && (
        (exe_valid && exe_is_load && exe_rf_we && (rf_raddr1 == exe_rf_waddr)) ||
        (mem_valid && mem_is_load && mem_rf_we && (rf_raddr1 == mem_rf_waddr))
    );
    wire rf_rdata2_hazard = use_rf_rdata2 && (
        (exe_valid && exe_is_load && exe_rf_we && (rf_raddr2 == exe_rf_waddr)) ||
        (mem_valid && mem_is_load && mem_rf_we && (rf_raddr2 == mem_rf_waddr))
    );

    assign id_ready_go = !rf_rdata1_hazard && !rf_rdata2_hazard;
    assign id_allow_in = !id_valid || id_ready_go && exe_allow_in;
    assign id_to_exe_valid = id_valid && id_ready_go;

    always @(posedge clk) begin
        if (reset) begin
            id_valid <= 1'b0;
            cancel_next <= 1'b0;
        end else if (br_cancel) begin
            id_valid <= 1'b0;
            cancel_next <= 1'b1;
        end else if (id_allow_in) begin
            id_valid <= if_to_id_valid;
        end
    end

    always @(posedge clk) begin
        if (id_allow_in && if_to_id_valid) begin
            id_reg <= if_to_id_bus;
            id_pred_br_taken <= if_to_id_bus[64];
            if (cancel_next) begin
                id_reg <= 0;
                cancel_next <= 0;
            end
        end else if (id_pred_br_taken) begin
            id_pred_br_taken <= 0;
        end
    end

    // BP Update
    assign upd_en = id_valid && id_ready_go && inst_is_br;
    assign upd_inst_addr = id_pc;
    assign upd_br_inst = inst_is_br;
    assign upd_cond_br_inst = inst_is_cond_br;
    assign upd_br_taken = br_taken;
    assign upd_br_target = br_target;

endmodule